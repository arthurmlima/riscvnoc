






out_W_controller_inst : entity work.out_W_controller
generic map(
    x_init      => x_init,
    y_init      => y_init,
    img_width   => img_width ,
    img_height  => img_height,
    n_frames    => n_frames  ,
    n_steps     => n_steps   ,
    pix_depth   => pix_depth
    )
port map(
	clk => clk,
	reset => reset,
	-- connections with the output controller
    oc_W_pixel   => W_input_CTRL_pixel  ,  
    oc_W_x_dest  => W_input_CTRL_x_dest ,  
    oc_W_y_dest  => W_input_CTRL_y_dest ,  
    oc_W_step    => W_input_CTRL_step   ,  
    oc_W_frame   => W_input_CTRL_frame  ,  
    oc_W_x_orig  => W_input_CTRL_x_orig ,  
    oc_W_y_orig  => W_input_CTRL_y_orig ,  
    oc_W_fb      => W_input_CTRL_fb     , 
     
    oc_W_new_msg => W_input_CTRL_req    ,  
    oc_W_ack     => W_input_CTRL_ack    ,
       
    -- connections to the next router
    i_W_pixel  => i_W_pixel,
    i_W_x_dest => i_W_x_dest,
    i_W_y_dest => i_W_y_dest,
    i_W_step   => i_W_step,
    i_W_frame  => i_W_frame,
    i_W_x_orig => i_W_x_orig,
    i_W_y_orig => i_W_y_orig,
    i_W_fb     => i_W_fb,
    i_W_req    => i_W_req,
    i_W_ack    => i_W_ack
    
);





























































































































































































































































































































































































































































































































































































































































































